connectix 